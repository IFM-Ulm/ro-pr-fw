`ifndef REPEAT_ASSIGN_OUTPUT_V
`define REPEAT_ASSIGN_OUTPUT_V 1

// Up to a number of 256 output ports, change only the following parameter. Otherwise extend the listing "_OUTPUT_REPEAT_..." as intended
`define MAX_PORTS_OUTPUT 32


`define SET_TEXT_OUTPUT(COUNTER) assign output_``COUNTER = w_output[COUNTER];

`define OUTPUT_REPEAT_ASSIGN(n) `_OUTPUT_REPEAT_``n
`define _OUTPUT_REPEAT_0
`define _OUTPUT_REPEAT_1  `SET_TEXT_OUTPUT(0)
`define _OUTPUT_REPEAT_2 `_OUTPUT_REPEAT_1 `SET_TEXT_OUTPUT(1)
`define _OUTPUT_REPEAT_3 `_OUTPUT_REPEAT_2 `SET_TEXT_OUTPUT(2)
`define _OUTPUT_REPEAT_4 `_OUTPUT_REPEAT_3 `SET_TEXT_OUTPUT(3)
`define _OUTPUT_REPEAT_5 `_OUTPUT_REPEAT_4 `SET_TEXT_OUTPUT(4)
`define _OUTPUT_REPEAT_6 `_OUTPUT_REPEAT_5 `SET_TEXT_OUTPUT(5)
`define _OUTPUT_REPEAT_7 `_OUTPUT_REPEAT_6 `SET_TEXT_OUTPUT(6)
`define _OUTPUT_REPEAT_8 `_OUTPUT_REPEAT_7 `SET_TEXT_OUTPUT(7)
`define _OUTPUT_REPEAT_9 `_OUTPUT_REPEAT_8 `SET_TEXT_OUTPUT(8)
`define _OUTPUT_REPEAT_10 `_OUTPUT_REPEAT_9 `SET_TEXT_OUTPUT(9)
`define _OUTPUT_REPEAT_11 `_OUTPUT_REPEAT_10 `SET_TEXT_OUTPUT(10)
`define _OUTPUT_REPEAT_12 `_OUTPUT_REPEAT_11 `SET_TEXT_OUTPUT(11)
`define _OUTPUT_REPEAT_13 `_OUTPUT_REPEAT_12 `SET_TEXT_OUTPUT(12)
`define _OUTPUT_REPEAT_14 `_OUTPUT_REPEAT_13 `SET_TEXT_OUTPUT(13)
`define _OUTPUT_REPEAT_15 `_OUTPUT_REPEAT_14 `SET_TEXT_OUTPUT(14)
`define _OUTPUT_REPEAT_16 `_OUTPUT_REPEAT_15 `SET_TEXT_OUTPUT(15)
`define _OUTPUT_REPEAT_17 `_OUTPUT_REPEAT_16 `SET_TEXT_OUTPUT(16)
`define _OUTPUT_REPEAT_18 `_OUTPUT_REPEAT_17 `SET_TEXT_OUTPUT(17)
`define _OUTPUT_REPEAT_19 `_OUTPUT_REPEAT_18 `SET_TEXT_OUTPUT(18)
`define _OUTPUT_REPEAT_20 `_OUTPUT_REPEAT_19 `SET_TEXT_OUTPUT(19)
`define _OUTPUT_REPEAT_21 `_OUTPUT_REPEAT_20 `SET_TEXT_OUTPUT(20)
`define _OUTPUT_REPEAT_22 `_OUTPUT_REPEAT_21 `SET_TEXT_OUTPUT(21)
`define _OUTPUT_REPEAT_23 `_OUTPUT_REPEAT_22 `SET_TEXT_OUTPUT(22)
`define _OUTPUT_REPEAT_24 `_OUTPUT_REPEAT_23 `SET_TEXT_OUTPUT(23)
`define _OUTPUT_REPEAT_25 `_OUTPUT_REPEAT_24 `SET_TEXT_OUTPUT(24)
`define _OUTPUT_REPEAT_26 `_OUTPUT_REPEAT_25 `SET_TEXT_OUTPUT(25)
`define _OUTPUT_REPEAT_27 `_OUTPUT_REPEAT_26 `SET_TEXT_OUTPUT(26)
`define _OUTPUT_REPEAT_28 `_OUTPUT_REPEAT_27 `SET_TEXT_OUTPUT(27)
`define _OUTPUT_REPEAT_29 `_OUTPUT_REPEAT_28 `SET_TEXT_OUTPUT(28)
`define _OUTPUT_REPEAT_30 `_OUTPUT_REPEAT_29 `SET_TEXT_OUTPUT(29)
`define _OUTPUT_REPEAT_31 `_OUTPUT_REPEAT_30 `SET_TEXT_OUTPUT(30)
`define _OUTPUT_REPEAT_32 `_OUTPUT_REPEAT_31 `SET_TEXT_OUTPUT(31)
`define _OUTPUT_REPEAT_33 `_OUTPUT_REPEAT_32 `SET_TEXT_OUTPUT(32)
`define _OUTPUT_REPEAT_34 `_OUTPUT_REPEAT_33 `SET_TEXT_OUTPUT(33)
`define _OUTPUT_REPEAT_35 `_OUTPUT_REPEAT_34 `SET_TEXT_OUTPUT(34)
`define _OUTPUT_REPEAT_36 `_OUTPUT_REPEAT_35 `SET_TEXT_OUTPUT(35)
`define _OUTPUT_REPEAT_37 `_OUTPUT_REPEAT_36 `SET_TEXT_OUTPUT(36)
`define _OUTPUT_REPEAT_38 `_OUTPUT_REPEAT_37 `SET_TEXT_OUTPUT(37)
`define _OUTPUT_REPEAT_39 `_OUTPUT_REPEAT_38 `SET_TEXT_OUTPUT(38)
`define _OUTPUT_REPEAT_40 `_OUTPUT_REPEAT_39 `SET_TEXT_OUTPUT(39)
`define _OUTPUT_REPEAT_41 `_OUTPUT_REPEAT_40 `SET_TEXT_OUTPUT(40)
`define _OUTPUT_REPEAT_42 `_OUTPUT_REPEAT_41 `SET_TEXT_OUTPUT(41)
`define _OUTPUT_REPEAT_43 `_OUTPUT_REPEAT_42 `SET_TEXT_OUTPUT(42)
`define _OUTPUT_REPEAT_44 `_OUTPUT_REPEAT_43 `SET_TEXT_OUTPUT(43)
`define _OUTPUT_REPEAT_45 `_OUTPUT_REPEAT_44 `SET_TEXT_OUTPUT(44)
`define _OUTPUT_REPEAT_46 `_OUTPUT_REPEAT_45 `SET_TEXT_OUTPUT(45)
`define _OUTPUT_REPEAT_47 `_OUTPUT_REPEAT_46 `SET_TEXT_OUTPUT(46)
`define _OUTPUT_REPEAT_48 `_OUTPUT_REPEAT_47 `SET_TEXT_OUTPUT(47)
`define _OUTPUT_REPEAT_49 `_OUTPUT_REPEAT_48 `SET_TEXT_OUTPUT(48)
`define _OUTPUT_REPEAT_50 `_OUTPUT_REPEAT_49 `SET_TEXT_OUTPUT(49)
`define _OUTPUT_REPEAT_51 `_OUTPUT_REPEAT_50 `SET_TEXT_OUTPUT(50)
`define _OUTPUT_REPEAT_52 `_OUTPUT_REPEAT_51 `SET_TEXT_OUTPUT(51)
`define _OUTPUT_REPEAT_53 `_OUTPUT_REPEAT_52 `SET_TEXT_OUTPUT(52)
`define _OUTPUT_REPEAT_54 `_OUTPUT_REPEAT_53 `SET_TEXT_OUTPUT(53)
`define _OUTPUT_REPEAT_55 `_OUTPUT_REPEAT_54 `SET_TEXT_OUTPUT(54)
`define _OUTPUT_REPEAT_56 `_OUTPUT_REPEAT_55 `SET_TEXT_OUTPUT(55)
`define _OUTPUT_REPEAT_57 `_OUTPUT_REPEAT_56 `SET_TEXT_OUTPUT(56)
`define _OUTPUT_REPEAT_58 `_OUTPUT_REPEAT_57 `SET_TEXT_OUTPUT(57)
`define _OUTPUT_REPEAT_59 `_OUTPUT_REPEAT_58 `SET_TEXT_OUTPUT(58)
`define _OUTPUT_REPEAT_60 `_OUTPUT_REPEAT_59 `SET_TEXT_OUTPUT(59)
`define _OUTPUT_REPEAT_61 `_OUTPUT_REPEAT_60 `SET_TEXT_OUTPUT(60)
`define _OUTPUT_REPEAT_62 `_OUTPUT_REPEAT_61 `SET_TEXT_OUTPUT(61)
`define _OUTPUT_REPEAT_63 `_OUTPUT_REPEAT_62 `SET_TEXT_OUTPUT(62)
`define _OUTPUT_REPEAT_64 `_OUTPUT_REPEAT_63 `SET_TEXT_OUTPUT(63)
`define _OUTPUT_REPEAT_65 `_OUTPUT_REPEAT_64 `SET_TEXT_OUTPUT(64)
`define _OUTPUT_REPEAT_66 `_OUTPUT_REPEAT_65 `SET_TEXT_OUTPUT(65)
`define _OUTPUT_REPEAT_67 `_OUTPUT_REPEAT_66 `SET_TEXT_OUTPUT(66)
`define _OUTPUT_REPEAT_68 `_OUTPUT_REPEAT_67 `SET_TEXT_OUTPUT(67)
`define _OUTPUT_REPEAT_69 `_OUTPUT_REPEAT_68 `SET_TEXT_OUTPUT(68)
`define _OUTPUT_REPEAT_70 `_OUTPUT_REPEAT_69 `SET_TEXT_OUTPUT(69)
`define _OUTPUT_REPEAT_71 `_OUTPUT_REPEAT_70 `SET_TEXT_OUTPUT(70)
`define _OUTPUT_REPEAT_72 `_OUTPUT_REPEAT_71 `SET_TEXT_OUTPUT(71)
`define _OUTPUT_REPEAT_73 `_OUTPUT_REPEAT_72 `SET_TEXT_OUTPUT(72)
`define _OUTPUT_REPEAT_74 `_OUTPUT_REPEAT_73 `SET_TEXT_OUTPUT(73)
`define _OUTPUT_REPEAT_75 `_OUTPUT_REPEAT_74 `SET_TEXT_OUTPUT(74)
`define _OUTPUT_REPEAT_76 `_OUTPUT_REPEAT_75 `SET_TEXT_OUTPUT(75)
`define _OUTPUT_REPEAT_77 `_OUTPUT_REPEAT_76 `SET_TEXT_OUTPUT(76)
`define _OUTPUT_REPEAT_78 `_OUTPUT_REPEAT_77 `SET_TEXT_OUTPUT(77)
`define _OUTPUT_REPEAT_79 `_OUTPUT_REPEAT_78 `SET_TEXT_OUTPUT(78)
`define _OUTPUT_REPEAT_80 `_OUTPUT_REPEAT_79 `SET_TEXT_OUTPUT(79)
`define _OUTPUT_REPEAT_81 `_OUTPUT_REPEAT_80 `SET_TEXT_OUTPUT(80)
`define _OUTPUT_REPEAT_82 `_OUTPUT_REPEAT_81 `SET_TEXT_OUTPUT(81)
`define _OUTPUT_REPEAT_83 `_OUTPUT_REPEAT_82 `SET_TEXT_OUTPUT(82)
`define _OUTPUT_REPEAT_84 `_OUTPUT_REPEAT_83 `SET_TEXT_OUTPUT(83)
`define _OUTPUT_REPEAT_85 `_OUTPUT_REPEAT_84 `SET_TEXT_OUTPUT(84)
`define _OUTPUT_REPEAT_86 `_OUTPUT_REPEAT_85 `SET_TEXT_OUTPUT(85)
`define _OUTPUT_REPEAT_87 `_OUTPUT_REPEAT_86 `SET_TEXT_OUTPUT(86)
`define _OUTPUT_REPEAT_88 `_OUTPUT_REPEAT_87 `SET_TEXT_OUTPUT(87)
`define _OUTPUT_REPEAT_89 `_OUTPUT_REPEAT_88 `SET_TEXT_OUTPUT(88)
`define _OUTPUT_REPEAT_90 `_OUTPUT_REPEAT_89 `SET_TEXT_OUTPUT(89)
`define _OUTPUT_REPEAT_91 `_OUTPUT_REPEAT_90 `SET_TEXT_OUTPUT(90)
`define _OUTPUT_REPEAT_92 `_OUTPUT_REPEAT_91 `SET_TEXT_OUTPUT(91)
`define _OUTPUT_REPEAT_93 `_OUTPUT_REPEAT_92 `SET_TEXT_OUTPUT(92)
`define _OUTPUT_REPEAT_94 `_OUTPUT_REPEAT_93 `SET_TEXT_OUTPUT(93)
`define _OUTPUT_REPEAT_95 `_OUTPUT_REPEAT_94 `SET_TEXT_OUTPUT(94)
`define _OUTPUT_REPEAT_96 `_OUTPUT_REPEAT_95 `SET_TEXT_OUTPUT(95)
`define _OUTPUT_REPEAT_97 `_OUTPUT_REPEAT_96 `SET_TEXT_OUTPUT(96)
`define _OUTPUT_REPEAT_98 `_OUTPUT_REPEAT_97 `SET_TEXT_OUTPUT(97)
`define _OUTPUT_REPEAT_99 `_OUTPUT_REPEAT_98 `SET_TEXT_OUTPUT(98)
`define _OUTPUT_REPEAT_100 `_OUTPUT_REPEAT_99 `SET_TEXT_OUTPUT(99)
`define _OUTPUT_REPEAT_101 `_OUTPUT_REPEAT_100 `SET_TEXT_OUTPUT(100)
`define _OUTPUT_REPEAT_102 `_OUTPUT_REPEAT_101 `SET_TEXT_OUTPUT(101)
`define _OUTPUT_REPEAT_103 `_OUTPUT_REPEAT_102 `SET_TEXT_OUTPUT(102)
`define _OUTPUT_REPEAT_104 `_OUTPUT_REPEAT_103 `SET_TEXT_OUTPUT(103)
`define _OUTPUT_REPEAT_105 `_OUTPUT_REPEAT_104 `SET_TEXT_OUTPUT(104)
`define _OUTPUT_REPEAT_106 `_OUTPUT_REPEAT_105 `SET_TEXT_OUTPUT(105)
`define _OUTPUT_REPEAT_107 `_OUTPUT_REPEAT_106 `SET_TEXT_OUTPUT(106)
`define _OUTPUT_REPEAT_108 `_OUTPUT_REPEAT_107 `SET_TEXT_OUTPUT(107)
`define _OUTPUT_REPEAT_109 `_OUTPUT_REPEAT_108 `SET_TEXT_OUTPUT(108)
`define _OUTPUT_REPEAT_110 `_OUTPUT_REPEAT_109 `SET_TEXT_OUTPUT(109)
`define _OUTPUT_REPEAT_111 `_OUTPUT_REPEAT_110 `SET_TEXT_OUTPUT(110)
`define _OUTPUT_REPEAT_112 `_OUTPUT_REPEAT_111 `SET_TEXT_OUTPUT(111)
`define _OUTPUT_REPEAT_113 `_OUTPUT_REPEAT_112 `SET_TEXT_OUTPUT(112)
`define _OUTPUT_REPEAT_114 `_OUTPUT_REPEAT_113 `SET_TEXT_OUTPUT(113)
`define _OUTPUT_REPEAT_115 `_OUTPUT_REPEAT_114 `SET_TEXT_OUTPUT(114)
`define _OUTPUT_REPEAT_116 `_OUTPUT_REPEAT_115 `SET_TEXT_OUTPUT(115)
`define _OUTPUT_REPEAT_117 `_OUTPUT_REPEAT_116 `SET_TEXT_OUTPUT(116)
`define _OUTPUT_REPEAT_118 `_OUTPUT_REPEAT_117 `SET_TEXT_OUTPUT(117)
`define _OUTPUT_REPEAT_119 `_OUTPUT_REPEAT_118 `SET_TEXT_OUTPUT(118)
`define _OUTPUT_REPEAT_120 `_OUTPUT_REPEAT_119 `SET_TEXT_OUTPUT(119)
`define _OUTPUT_REPEAT_121 `_OUTPUT_REPEAT_120 `SET_TEXT_OUTPUT(120)
`define _OUTPUT_REPEAT_122 `_OUTPUT_REPEAT_121 `SET_TEXT_OUTPUT(121)
`define _OUTPUT_REPEAT_123 `_OUTPUT_REPEAT_122 `SET_TEXT_OUTPUT(122)
`define _OUTPUT_REPEAT_124 `_OUTPUT_REPEAT_123 `SET_TEXT_OUTPUT(123)
`define _OUTPUT_REPEAT_125 `_OUTPUT_REPEAT_124 `SET_TEXT_OUTPUT(124)
`define _OUTPUT_REPEAT_126 `_OUTPUT_REPEAT_125 `SET_TEXT_OUTPUT(125)
`define _OUTPUT_REPEAT_127 `_OUTPUT_REPEAT_126 `SET_TEXT_OUTPUT(126)
`define _OUTPUT_REPEAT_128 `_OUTPUT_REPEAT_127 `SET_TEXT_OUTPUT(127)
`define _OUTPUT_REPEAT_129 `_OUTPUT_REPEAT_128 `SET_TEXT_OUTPUT(128)
`define _OUTPUT_REPEAT_130 `_OUTPUT_REPEAT_129 `SET_TEXT_OUTPUT(129)
`define _OUTPUT_REPEAT_131 `_OUTPUT_REPEAT_130 `SET_TEXT_OUTPUT(130)
`define _OUTPUT_REPEAT_132 `_OUTPUT_REPEAT_131 `SET_TEXT_OUTPUT(131)
`define _OUTPUT_REPEAT_133 `_OUTPUT_REPEAT_132 `SET_TEXT_OUTPUT(132)
`define _OUTPUT_REPEAT_134 `_OUTPUT_REPEAT_133 `SET_TEXT_OUTPUT(133)
`define _OUTPUT_REPEAT_135 `_OUTPUT_REPEAT_134 `SET_TEXT_OUTPUT(134)
`define _OUTPUT_REPEAT_136 `_OUTPUT_REPEAT_135 `SET_TEXT_OUTPUT(135)
`define _OUTPUT_REPEAT_137 `_OUTPUT_REPEAT_136 `SET_TEXT_OUTPUT(136)
`define _OUTPUT_REPEAT_138 `_OUTPUT_REPEAT_137 `SET_TEXT_OUTPUT(137)
`define _OUTPUT_REPEAT_139 `_OUTPUT_REPEAT_138 `SET_TEXT_OUTPUT(138)
`define _OUTPUT_REPEAT_140 `_OUTPUT_REPEAT_139 `SET_TEXT_OUTPUT(139)
`define _OUTPUT_REPEAT_141 `_OUTPUT_REPEAT_140 `SET_TEXT_OUTPUT(140)
`define _OUTPUT_REPEAT_142 `_OUTPUT_REPEAT_141 `SET_TEXT_OUTPUT(141)
`define _OUTPUT_REPEAT_143 `_OUTPUT_REPEAT_142 `SET_TEXT_OUTPUT(142)
`define _OUTPUT_REPEAT_144 `_OUTPUT_REPEAT_143 `SET_TEXT_OUTPUT(143)
`define _OUTPUT_REPEAT_145 `_OUTPUT_REPEAT_144 `SET_TEXT_OUTPUT(144)
`define _OUTPUT_REPEAT_146 `_OUTPUT_REPEAT_145 `SET_TEXT_OUTPUT(145)
`define _OUTPUT_REPEAT_147 `_OUTPUT_REPEAT_146 `SET_TEXT_OUTPUT(146)
`define _OUTPUT_REPEAT_148 `_OUTPUT_REPEAT_147 `SET_TEXT_OUTPUT(147)
`define _OUTPUT_REPEAT_149 `_OUTPUT_REPEAT_148 `SET_TEXT_OUTPUT(148)
`define _OUTPUT_REPEAT_150 `_OUTPUT_REPEAT_149 `SET_TEXT_OUTPUT(149)
`define _OUTPUT_REPEAT_151 `_OUTPUT_REPEAT_150 `SET_TEXT_OUTPUT(150)
`define _OUTPUT_REPEAT_152 `_OUTPUT_REPEAT_151 `SET_TEXT_OUTPUT(151)
`define _OUTPUT_REPEAT_153 `_OUTPUT_REPEAT_152 `SET_TEXT_OUTPUT(152)
`define _OUTPUT_REPEAT_154 `_OUTPUT_REPEAT_153 `SET_TEXT_OUTPUT(153)
`define _OUTPUT_REPEAT_155 `_OUTPUT_REPEAT_154 `SET_TEXT_OUTPUT(154)
`define _OUTPUT_REPEAT_156 `_OUTPUT_REPEAT_155 `SET_TEXT_OUTPUT(155)
`define _OUTPUT_REPEAT_157 `_OUTPUT_REPEAT_156 `SET_TEXT_OUTPUT(156)
`define _OUTPUT_REPEAT_158 `_OUTPUT_REPEAT_157 `SET_TEXT_OUTPUT(157)
`define _OUTPUT_REPEAT_159 `_OUTPUT_REPEAT_158 `SET_TEXT_OUTPUT(158)
`define _OUTPUT_REPEAT_160 `_OUTPUT_REPEAT_159 `SET_TEXT_OUTPUT(159)
`define _OUTPUT_REPEAT_161 `_OUTPUT_REPEAT_160 `SET_TEXT_OUTPUT(160)
`define _OUTPUT_REPEAT_162 `_OUTPUT_REPEAT_161 `SET_TEXT_OUTPUT(161)
`define _OUTPUT_REPEAT_163 `_OUTPUT_REPEAT_162 `SET_TEXT_OUTPUT(162)
`define _OUTPUT_REPEAT_164 `_OUTPUT_REPEAT_163 `SET_TEXT_OUTPUT(163)
`define _OUTPUT_REPEAT_165 `_OUTPUT_REPEAT_164 `SET_TEXT_OUTPUT(164)
`define _OUTPUT_REPEAT_166 `_OUTPUT_REPEAT_165 `SET_TEXT_OUTPUT(165)
`define _OUTPUT_REPEAT_167 `_OUTPUT_REPEAT_166 `SET_TEXT_OUTPUT(166)
`define _OUTPUT_REPEAT_168 `_OUTPUT_REPEAT_167 `SET_TEXT_OUTPUT(167)
`define _OUTPUT_REPEAT_169 `_OUTPUT_REPEAT_168 `SET_TEXT_OUTPUT(168)
`define _OUTPUT_REPEAT_170 `_OUTPUT_REPEAT_169 `SET_TEXT_OUTPUT(169)
`define _OUTPUT_REPEAT_171 `_OUTPUT_REPEAT_170 `SET_TEXT_OUTPUT(170)
`define _OUTPUT_REPEAT_172 `_OUTPUT_REPEAT_171 `SET_TEXT_OUTPUT(171)
`define _OUTPUT_REPEAT_173 `_OUTPUT_REPEAT_172 `SET_TEXT_OUTPUT(172)
`define _OUTPUT_REPEAT_174 `_OUTPUT_REPEAT_173 `SET_TEXT_OUTPUT(173)
`define _OUTPUT_REPEAT_175 `_OUTPUT_REPEAT_174 `SET_TEXT_OUTPUT(174)
`define _OUTPUT_REPEAT_176 `_OUTPUT_REPEAT_175 `SET_TEXT_OUTPUT(175)
`define _OUTPUT_REPEAT_177 `_OUTPUT_REPEAT_176 `SET_TEXT_OUTPUT(176)
`define _OUTPUT_REPEAT_178 `_OUTPUT_REPEAT_177 `SET_TEXT_OUTPUT(177)
`define _OUTPUT_REPEAT_179 `_OUTPUT_REPEAT_178 `SET_TEXT_OUTPUT(178)
`define _OUTPUT_REPEAT_180 `_OUTPUT_REPEAT_179 `SET_TEXT_OUTPUT(179)
`define _OUTPUT_REPEAT_181 `_OUTPUT_REPEAT_180 `SET_TEXT_OUTPUT(180)
`define _OUTPUT_REPEAT_182 `_OUTPUT_REPEAT_181 `SET_TEXT_OUTPUT(181)
`define _OUTPUT_REPEAT_183 `_OUTPUT_REPEAT_182 `SET_TEXT_OUTPUT(182)
`define _OUTPUT_REPEAT_184 `_OUTPUT_REPEAT_183 `SET_TEXT_OUTPUT(183)
`define _OUTPUT_REPEAT_185 `_OUTPUT_REPEAT_184 `SET_TEXT_OUTPUT(184)
`define _OUTPUT_REPEAT_186 `_OUTPUT_REPEAT_185 `SET_TEXT_OUTPUT(185)
`define _OUTPUT_REPEAT_187 `_OUTPUT_REPEAT_186 `SET_TEXT_OUTPUT(186)
`define _OUTPUT_REPEAT_188 `_OUTPUT_REPEAT_187 `SET_TEXT_OUTPUT(187)
`define _OUTPUT_REPEAT_189 `_OUTPUT_REPEAT_188 `SET_TEXT_OUTPUT(188)
`define _OUTPUT_REPEAT_190 `_OUTPUT_REPEAT_189 `SET_TEXT_OUTPUT(189)
`define _OUTPUT_REPEAT_191 `_OUTPUT_REPEAT_190 `SET_TEXT_OUTPUT(190)
`define _OUTPUT_REPEAT_192 `_OUTPUT_REPEAT_191 `SET_TEXT_OUTPUT(191)
`define _OUTPUT_REPEAT_193 `_OUTPUT_REPEAT_192 `SET_TEXT_OUTPUT(192)
`define _OUTPUT_REPEAT_194 `_OUTPUT_REPEAT_193 `SET_TEXT_OUTPUT(193)
`define _OUTPUT_REPEAT_195 `_OUTPUT_REPEAT_194 `SET_TEXT_OUTPUT(194)
`define _OUTPUT_REPEAT_196 `_OUTPUT_REPEAT_195 `SET_TEXT_OUTPUT(195)
`define _OUTPUT_REPEAT_197 `_OUTPUT_REPEAT_196 `SET_TEXT_OUTPUT(196)
`define _OUTPUT_REPEAT_198 `_OUTPUT_REPEAT_197 `SET_TEXT_OUTPUT(197)
`define _OUTPUT_REPEAT_199 `_OUTPUT_REPEAT_198 `SET_TEXT_OUTPUT(198)
`define _OUTPUT_REPEAT_200 `_OUTPUT_REPEAT_199 `SET_TEXT_OUTPUT(199)
`define _OUTPUT_REPEAT_201 `_OUTPUT_REPEAT_200 `SET_TEXT_OUTPUT(200)
`define _OUTPUT_REPEAT_202 `_OUTPUT_REPEAT_201 `SET_TEXT_OUTPUT(201)
`define _OUTPUT_REPEAT_203 `_OUTPUT_REPEAT_202 `SET_TEXT_OUTPUT(202)
`define _OUTPUT_REPEAT_204 `_OUTPUT_REPEAT_203 `SET_TEXT_OUTPUT(203)
`define _OUTPUT_REPEAT_205 `_OUTPUT_REPEAT_204 `SET_TEXT_OUTPUT(204)
`define _OUTPUT_REPEAT_206 `_OUTPUT_REPEAT_205 `SET_TEXT_OUTPUT(205)
`define _OUTPUT_REPEAT_207 `_OUTPUT_REPEAT_206 `SET_TEXT_OUTPUT(206)
`define _OUTPUT_REPEAT_208 `_OUTPUT_REPEAT_207 `SET_TEXT_OUTPUT(207)
`define _OUTPUT_REPEAT_209 `_OUTPUT_REPEAT_208 `SET_TEXT_OUTPUT(208)
`define _OUTPUT_REPEAT_210 `_OUTPUT_REPEAT_209 `SET_TEXT_OUTPUT(209)
`define _OUTPUT_REPEAT_211 `_OUTPUT_REPEAT_210 `SET_TEXT_OUTPUT(210)
`define _OUTPUT_REPEAT_212 `_OUTPUT_REPEAT_211 `SET_TEXT_OUTPUT(211)
`define _OUTPUT_REPEAT_213 `_OUTPUT_REPEAT_212 `SET_TEXT_OUTPUT(212)
`define _OUTPUT_REPEAT_214 `_OUTPUT_REPEAT_213 `SET_TEXT_OUTPUT(213)
`define _OUTPUT_REPEAT_215 `_OUTPUT_REPEAT_214 `SET_TEXT_OUTPUT(214)
`define _OUTPUT_REPEAT_216 `_OUTPUT_REPEAT_215 `SET_TEXT_OUTPUT(215)
`define _OUTPUT_REPEAT_217 `_OUTPUT_REPEAT_216 `SET_TEXT_OUTPUT(216)
`define _OUTPUT_REPEAT_218 `_OUTPUT_REPEAT_217 `SET_TEXT_OUTPUT(217)
`define _OUTPUT_REPEAT_219 `_OUTPUT_REPEAT_218 `SET_TEXT_OUTPUT(218)
`define _OUTPUT_REPEAT_220 `_OUTPUT_REPEAT_219 `SET_TEXT_OUTPUT(219)
`define _OUTPUT_REPEAT_221 `_OUTPUT_REPEAT_220 `SET_TEXT_OUTPUT(220)
`define _OUTPUT_REPEAT_222 `_OUTPUT_REPEAT_221 `SET_TEXT_OUTPUT(221)
`define _OUTPUT_REPEAT_223 `_OUTPUT_REPEAT_222 `SET_TEXT_OUTPUT(222)
`define _OUTPUT_REPEAT_224 `_OUTPUT_REPEAT_223 `SET_TEXT_OUTPUT(223)
`define _OUTPUT_REPEAT_225 `_OUTPUT_REPEAT_224 `SET_TEXT_OUTPUT(224)
`define _OUTPUT_REPEAT_226 `_OUTPUT_REPEAT_225 `SET_TEXT_OUTPUT(225)
`define _OUTPUT_REPEAT_227 `_OUTPUT_REPEAT_226 `SET_TEXT_OUTPUT(226)
`define _OUTPUT_REPEAT_228 `_OUTPUT_REPEAT_227 `SET_TEXT_OUTPUT(227)
`define _OUTPUT_REPEAT_229 `_OUTPUT_REPEAT_228 `SET_TEXT_OUTPUT(228)
`define _OUTPUT_REPEAT_230 `_OUTPUT_REPEAT_229 `SET_TEXT_OUTPUT(229)
`define _OUTPUT_REPEAT_231 `_OUTPUT_REPEAT_230 `SET_TEXT_OUTPUT(230)
`define _OUTPUT_REPEAT_232 `_OUTPUT_REPEAT_231 `SET_TEXT_OUTPUT(231)
`define _OUTPUT_REPEAT_233 `_OUTPUT_REPEAT_232 `SET_TEXT_OUTPUT(232)
`define _OUTPUT_REPEAT_234 `_OUTPUT_REPEAT_233 `SET_TEXT_OUTPUT(233)
`define _OUTPUT_REPEAT_235 `_OUTPUT_REPEAT_234 `SET_TEXT_OUTPUT(234)
`define _OUTPUT_REPEAT_236 `_OUTPUT_REPEAT_235 `SET_TEXT_OUTPUT(235)
`define _OUTPUT_REPEAT_237 `_OUTPUT_REPEAT_236 `SET_TEXT_OUTPUT(236)
`define _OUTPUT_REPEAT_238 `_OUTPUT_REPEAT_237 `SET_TEXT_OUTPUT(237)
`define _OUTPUT_REPEAT_239 `_OUTPUT_REPEAT_238 `SET_TEXT_OUTPUT(238)
`define _OUTPUT_REPEAT_240 `_OUTPUT_REPEAT_239 `SET_TEXT_OUTPUT(239)
`define _OUTPUT_REPEAT_241 `_OUTPUT_REPEAT_240 `SET_TEXT_OUTPUT(240)
`define _OUTPUT_REPEAT_242 `_OUTPUT_REPEAT_241 `SET_TEXT_OUTPUT(241)
`define _OUTPUT_REPEAT_243 `_OUTPUT_REPEAT_242 `SET_TEXT_OUTPUT(242)
`define _OUTPUT_REPEAT_244 `_OUTPUT_REPEAT_243 `SET_TEXT_OUTPUT(243)
`define _OUTPUT_REPEAT_245 `_OUTPUT_REPEAT_244 `SET_TEXT_OUTPUT(244)
`define _OUTPUT_REPEAT_246 `_OUTPUT_REPEAT_245 `SET_TEXT_OUTPUT(245)
`define _OUTPUT_REPEAT_247 `_OUTPUT_REPEAT_246 `SET_TEXT_OUTPUT(246)
`define _OUTPUT_REPEAT_248 `_OUTPUT_REPEAT_247 `SET_TEXT_OUTPUT(247)
`define _OUTPUT_REPEAT_249 `_OUTPUT_REPEAT_248 `SET_TEXT_OUTPUT(248)
`define _OUTPUT_REPEAT_250 `_OUTPUT_REPEAT_249 `SET_TEXT_OUTPUT(249)
`define _OUTPUT_REPEAT_251 `_OUTPUT_REPEAT_250 `SET_TEXT_OUTPUT(250)
`define _OUTPUT_REPEAT_252 `_OUTPUT_REPEAT_251 `SET_TEXT_OUTPUT(251)
`define _OUTPUT_REPEAT_253 `_OUTPUT_REPEAT_252 `SET_TEXT_OUTPUT(252)
`define _OUTPUT_REPEAT_254 `_OUTPUT_REPEAT_253 `SET_TEXT_OUTPUT(253)
`define _OUTPUT_REPEAT_255 `_OUTPUT_REPEAT_254 `SET_TEXT_OUTPUT(254)
`define _OUTPUT_REPEAT_256 `_OUTPUT_REPEAT_255 `SET_TEXT_OUTPUT(255)


`endif