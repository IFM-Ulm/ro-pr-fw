module PR_empty (
		input wire [31:0] counting,
		output wire [31:0] RO_out
);

assign RO_out = 0;

endmodule