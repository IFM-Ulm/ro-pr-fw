`ifndef REPEAT_ASSIGN_INPUT_V
`define REPEAT_ASSIGN_INPUT_V 1

// Up to a number of 256 input ports, change only the following parameter. Otherwise extend the listing "_INPUT_REPEAT_..." as intended
`define MAX_PORTS_INPUT 32


`define SET_TEXT_INPUT(COUNTER) assign w_input[COUNTER] = input_``COUNTER;

`define INPUT_REPEAT_ASSIGN(n) `_INPUT_REPEAT_``n
`define _INPUT_REPEAT_0
`define _INPUT_REPEAT_1  `SET_TEXT_INPUT(0)
`define _INPUT_REPEAT_2 `_INPUT_REPEAT_1 `SET_TEXT_INPUT(1)
`define _INPUT_REPEAT_3 `_INPUT_REPEAT_2 `SET_TEXT_INPUT(2)
`define _INPUT_REPEAT_4 `_INPUT_REPEAT_3 `SET_TEXT_INPUT(3)
`define _INPUT_REPEAT_5 `_INPUT_REPEAT_4 `SET_TEXT_INPUT(4)
`define _INPUT_REPEAT_6 `_INPUT_REPEAT_5 `SET_TEXT_INPUT(5)
`define _INPUT_REPEAT_7 `_INPUT_REPEAT_6 `SET_TEXT_INPUT(6)
`define _INPUT_REPEAT_8 `_INPUT_REPEAT_7 `SET_TEXT_INPUT(7)
`define _INPUT_REPEAT_9 `_INPUT_REPEAT_8 `SET_TEXT_INPUT(8)
`define _INPUT_REPEAT_10 `_INPUT_REPEAT_9 `SET_TEXT_INPUT(9)
`define _INPUT_REPEAT_11 `_INPUT_REPEAT_10 `SET_TEXT_INPUT(10)
`define _INPUT_REPEAT_12 `_INPUT_REPEAT_11 `SET_TEXT_INPUT(11)
`define _INPUT_REPEAT_13 `_INPUT_REPEAT_12 `SET_TEXT_INPUT(12)
`define _INPUT_REPEAT_14 `_INPUT_REPEAT_13 `SET_TEXT_INPUT(13)
`define _INPUT_REPEAT_15 `_INPUT_REPEAT_14 `SET_TEXT_INPUT(14)
`define _INPUT_REPEAT_16 `_INPUT_REPEAT_15 `SET_TEXT_INPUT(15)
`define _INPUT_REPEAT_17 `_INPUT_REPEAT_16 `SET_TEXT_INPUT(16)
`define _INPUT_REPEAT_18 `_INPUT_REPEAT_17 `SET_TEXT_INPUT(17)
`define _INPUT_REPEAT_19 `_INPUT_REPEAT_18 `SET_TEXT_INPUT(18)
`define _INPUT_REPEAT_20 `_INPUT_REPEAT_19 `SET_TEXT_INPUT(19)
`define _INPUT_REPEAT_21 `_INPUT_REPEAT_20 `SET_TEXT_INPUT(20)
`define _INPUT_REPEAT_22 `_INPUT_REPEAT_21 `SET_TEXT_INPUT(21)
`define _INPUT_REPEAT_23 `_INPUT_REPEAT_22 `SET_TEXT_INPUT(22)
`define _INPUT_REPEAT_24 `_INPUT_REPEAT_23 `SET_TEXT_INPUT(23)
`define _INPUT_REPEAT_25 `_INPUT_REPEAT_24 `SET_TEXT_INPUT(24)
`define _INPUT_REPEAT_26 `_INPUT_REPEAT_25 `SET_TEXT_INPUT(25)
`define _INPUT_REPEAT_27 `_INPUT_REPEAT_26 `SET_TEXT_INPUT(26)
`define _INPUT_REPEAT_28 `_INPUT_REPEAT_27 `SET_TEXT_INPUT(27)
`define _INPUT_REPEAT_29 `_INPUT_REPEAT_28 `SET_TEXT_INPUT(28)
`define _INPUT_REPEAT_30 `_INPUT_REPEAT_29 `SET_TEXT_INPUT(29)
`define _INPUT_REPEAT_31 `_INPUT_REPEAT_30 `SET_TEXT_INPUT(30)
`define _INPUT_REPEAT_32 `_INPUT_REPEAT_31 `SET_TEXT_INPUT(31)
`define _INPUT_REPEAT_33 `_INPUT_REPEAT_32 `SET_TEXT_INPUT(32)
`define _INPUT_REPEAT_34 `_INPUT_REPEAT_33 `SET_TEXT_INPUT(33)
`define _INPUT_REPEAT_35 `_INPUT_REPEAT_34 `SET_TEXT_INPUT(34)
`define _INPUT_REPEAT_36 `_INPUT_REPEAT_35 `SET_TEXT_INPUT(35)
`define _INPUT_REPEAT_37 `_INPUT_REPEAT_36 `SET_TEXT_INPUT(36)
`define _INPUT_REPEAT_38 `_INPUT_REPEAT_37 `SET_TEXT_INPUT(37)
`define _INPUT_REPEAT_39 `_INPUT_REPEAT_38 `SET_TEXT_INPUT(38)
`define _INPUT_REPEAT_40 `_INPUT_REPEAT_39 `SET_TEXT_INPUT(39)
`define _INPUT_REPEAT_41 `_INPUT_REPEAT_40 `SET_TEXT_INPUT(40)
`define _INPUT_REPEAT_42 `_INPUT_REPEAT_41 `SET_TEXT_INPUT(41)
`define _INPUT_REPEAT_43 `_INPUT_REPEAT_42 `SET_TEXT_INPUT(42)
`define _INPUT_REPEAT_44 `_INPUT_REPEAT_43 `SET_TEXT_INPUT(43)
`define _INPUT_REPEAT_45 `_INPUT_REPEAT_44 `SET_TEXT_INPUT(44)
`define _INPUT_REPEAT_46 `_INPUT_REPEAT_45 `SET_TEXT_INPUT(45)
`define _INPUT_REPEAT_47 `_INPUT_REPEAT_46 `SET_TEXT_INPUT(46)
`define _INPUT_REPEAT_48 `_INPUT_REPEAT_47 `SET_TEXT_INPUT(47)
`define _INPUT_REPEAT_49 `_INPUT_REPEAT_48 `SET_TEXT_INPUT(48)
`define _INPUT_REPEAT_50 `_INPUT_REPEAT_49 `SET_TEXT_INPUT(49)
`define _INPUT_REPEAT_51 `_INPUT_REPEAT_50 `SET_TEXT_INPUT(50)
`define _INPUT_REPEAT_52 `_INPUT_REPEAT_51 `SET_TEXT_INPUT(51)
`define _INPUT_REPEAT_53 `_INPUT_REPEAT_52 `SET_TEXT_INPUT(52)
`define _INPUT_REPEAT_54 `_INPUT_REPEAT_53 `SET_TEXT_INPUT(53)
`define _INPUT_REPEAT_55 `_INPUT_REPEAT_54 `SET_TEXT_INPUT(54)
`define _INPUT_REPEAT_56 `_INPUT_REPEAT_55 `SET_TEXT_INPUT(55)
`define _INPUT_REPEAT_57 `_INPUT_REPEAT_56 `SET_TEXT_INPUT(56)
`define _INPUT_REPEAT_58 `_INPUT_REPEAT_57 `SET_TEXT_INPUT(57)
`define _INPUT_REPEAT_59 `_INPUT_REPEAT_58 `SET_TEXT_INPUT(58)
`define _INPUT_REPEAT_60 `_INPUT_REPEAT_59 `SET_TEXT_INPUT(59)
`define _INPUT_REPEAT_61 `_INPUT_REPEAT_60 `SET_TEXT_INPUT(60)
`define _INPUT_REPEAT_62 `_INPUT_REPEAT_61 `SET_TEXT_INPUT(61)
`define _INPUT_REPEAT_63 `_INPUT_REPEAT_62 `SET_TEXT_INPUT(62)
`define _INPUT_REPEAT_64 `_INPUT_REPEAT_63 `SET_TEXT_INPUT(63)
`define _INPUT_REPEAT_65 `_INPUT_REPEAT_64 `SET_TEXT_INPUT(64)
`define _INPUT_REPEAT_66 `_INPUT_REPEAT_65 `SET_TEXT_INPUT(65)
`define _INPUT_REPEAT_67 `_INPUT_REPEAT_66 `SET_TEXT_INPUT(66)
`define _INPUT_REPEAT_68 `_INPUT_REPEAT_67 `SET_TEXT_INPUT(67)
`define _INPUT_REPEAT_69 `_INPUT_REPEAT_68 `SET_TEXT_INPUT(68)
`define _INPUT_REPEAT_70 `_INPUT_REPEAT_69 `SET_TEXT_INPUT(69)
`define _INPUT_REPEAT_71 `_INPUT_REPEAT_70 `SET_TEXT_INPUT(70)
`define _INPUT_REPEAT_72 `_INPUT_REPEAT_71 `SET_TEXT_INPUT(71)
`define _INPUT_REPEAT_73 `_INPUT_REPEAT_72 `SET_TEXT_INPUT(72)
`define _INPUT_REPEAT_74 `_INPUT_REPEAT_73 `SET_TEXT_INPUT(73)
`define _INPUT_REPEAT_75 `_INPUT_REPEAT_74 `SET_TEXT_INPUT(74)
`define _INPUT_REPEAT_76 `_INPUT_REPEAT_75 `SET_TEXT_INPUT(75)
`define _INPUT_REPEAT_77 `_INPUT_REPEAT_76 `SET_TEXT_INPUT(76)
`define _INPUT_REPEAT_78 `_INPUT_REPEAT_77 `SET_TEXT_INPUT(77)
`define _INPUT_REPEAT_79 `_INPUT_REPEAT_78 `SET_TEXT_INPUT(78)
`define _INPUT_REPEAT_80 `_INPUT_REPEAT_79 `SET_TEXT_INPUT(79)
`define _INPUT_REPEAT_81 `_INPUT_REPEAT_80 `SET_TEXT_INPUT(80)
`define _INPUT_REPEAT_82 `_INPUT_REPEAT_81 `SET_TEXT_INPUT(81)
`define _INPUT_REPEAT_83 `_INPUT_REPEAT_82 `SET_TEXT_INPUT(82)
`define _INPUT_REPEAT_84 `_INPUT_REPEAT_83 `SET_TEXT_INPUT(83)
`define _INPUT_REPEAT_85 `_INPUT_REPEAT_84 `SET_TEXT_INPUT(84)
`define _INPUT_REPEAT_86 `_INPUT_REPEAT_85 `SET_TEXT_INPUT(85)
`define _INPUT_REPEAT_87 `_INPUT_REPEAT_86 `SET_TEXT_INPUT(86)
`define _INPUT_REPEAT_88 `_INPUT_REPEAT_87 `SET_TEXT_INPUT(87)
`define _INPUT_REPEAT_89 `_INPUT_REPEAT_88 `SET_TEXT_INPUT(88)
`define _INPUT_REPEAT_90 `_INPUT_REPEAT_89 `SET_TEXT_INPUT(89)
`define _INPUT_REPEAT_91 `_INPUT_REPEAT_90 `SET_TEXT_INPUT(90)
`define _INPUT_REPEAT_92 `_INPUT_REPEAT_91 `SET_TEXT_INPUT(91)
`define _INPUT_REPEAT_93 `_INPUT_REPEAT_92 `SET_TEXT_INPUT(92)
`define _INPUT_REPEAT_94 `_INPUT_REPEAT_93 `SET_TEXT_INPUT(93)
`define _INPUT_REPEAT_95 `_INPUT_REPEAT_94 `SET_TEXT_INPUT(94)
`define _INPUT_REPEAT_96 `_INPUT_REPEAT_95 `SET_TEXT_INPUT(95)
`define _INPUT_REPEAT_97 `_INPUT_REPEAT_96 `SET_TEXT_INPUT(96)
`define _INPUT_REPEAT_98 `_INPUT_REPEAT_97 `SET_TEXT_INPUT(97)
`define _INPUT_REPEAT_99 `_INPUT_REPEAT_98 `SET_TEXT_INPUT(98)
`define _INPUT_REPEAT_100 `_INPUT_REPEAT_99 `SET_TEXT_INPUT(99)
`define _INPUT_REPEAT_101 `_INPUT_REPEAT_100 `SET_TEXT_INPUT(100)
`define _INPUT_REPEAT_102 `_INPUT_REPEAT_101 `SET_TEXT_INPUT(101)
`define _INPUT_REPEAT_103 `_INPUT_REPEAT_102 `SET_TEXT_INPUT(102)
`define _INPUT_REPEAT_104 `_INPUT_REPEAT_103 `SET_TEXT_INPUT(103)
`define _INPUT_REPEAT_105 `_INPUT_REPEAT_104 `SET_TEXT_INPUT(104)
`define _INPUT_REPEAT_106 `_INPUT_REPEAT_105 `SET_TEXT_INPUT(105)
`define _INPUT_REPEAT_107 `_INPUT_REPEAT_106 `SET_TEXT_INPUT(106)
`define _INPUT_REPEAT_108 `_INPUT_REPEAT_107 `SET_TEXT_INPUT(107)
`define _INPUT_REPEAT_109 `_INPUT_REPEAT_108 `SET_TEXT_INPUT(108)
`define _INPUT_REPEAT_110 `_INPUT_REPEAT_109 `SET_TEXT_INPUT(109)
`define _INPUT_REPEAT_111 `_INPUT_REPEAT_110 `SET_TEXT_INPUT(110)
`define _INPUT_REPEAT_112 `_INPUT_REPEAT_111 `SET_TEXT_INPUT(111)
`define _INPUT_REPEAT_113 `_INPUT_REPEAT_112 `SET_TEXT_INPUT(112)
`define _INPUT_REPEAT_114 `_INPUT_REPEAT_113 `SET_TEXT_INPUT(113)
`define _INPUT_REPEAT_115 `_INPUT_REPEAT_114 `SET_TEXT_INPUT(114)
`define _INPUT_REPEAT_116 `_INPUT_REPEAT_115 `SET_TEXT_INPUT(115)
`define _INPUT_REPEAT_117 `_INPUT_REPEAT_116 `SET_TEXT_INPUT(116)
`define _INPUT_REPEAT_118 `_INPUT_REPEAT_117 `SET_TEXT_INPUT(117)
`define _INPUT_REPEAT_119 `_INPUT_REPEAT_118 `SET_TEXT_INPUT(118)
`define _INPUT_REPEAT_120 `_INPUT_REPEAT_119 `SET_TEXT_INPUT(119)
`define _INPUT_REPEAT_121 `_INPUT_REPEAT_120 `SET_TEXT_INPUT(120)
`define _INPUT_REPEAT_122 `_INPUT_REPEAT_121 `SET_TEXT_INPUT(121)
`define _INPUT_REPEAT_123 `_INPUT_REPEAT_122 `SET_TEXT_INPUT(122)
`define _INPUT_REPEAT_124 `_INPUT_REPEAT_123 `SET_TEXT_INPUT(123)
`define _INPUT_REPEAT_125 `_INPUT_REPEAT_124 `SET_TEXT_INPUT(124)
`define _INPUT_REPEAT_126 `_INPUT_REPEAT_125 `SET_TEXT_INPUT(125)
`define _INPUT_REPEAT_127 `_INPUT_REPEAT_126 `SET_TEXT_INPUT(126)
`define _INPUT_REPEAT_128 `_INPUT_REPEAT_127 `SET_TEXT_INPUT(127)
`define _INPUT_REPEAT_129 `_INPUT_REPEAT_128 `SET_TEXT_INPUT(128)
`define _INPUT_REPEAT_130 `_INPUT_REPEAT_129 `SET_TEXT_INPUT(129)
`define _INPUT_REPEAT_131 `_INPUT_REPEAT_130 `SET_TEXT_INPUT(130)
`define _INPUT_REPEAT_132 `_INPUT_REPEAT_131 `SET_TEXT_INPUT(131)
`define _INPUT_REPEAT_133 `_INPUT_REPEAT_132 `SET_TEXT_INPUT(132)
`define _INPUT_REPEAT_134 `_INPUT_REPEAT_133 `SET_TEXT_INPUT(133)
`define _INPUT_REPEAT_135 `_INPUT_REPEAT_134 `SET_TEXT_INPUT(134)
`define _INPUT_REPEAT_136 `_INPUT_REPEAT_135 `SET_TEXT_INPUT(135)
`define _INPUT_REPEAT_137 `_INPUT_REPEAT_136 `SET_TEXT_INPUT(136)
`define _INPUT_REPEAT_138 `_INPUT_REPEAT_137 `SET_TEXT_INPUT(137)
`define _INPUT_REPEAT_139 `_INPUT_REPEAT_138 `SET_TEXT_INPUT(138)
`define _INPUT_REPEAT_140 `_INPUT_REPEAT_139 `SET_TEXT_INPUT(139)
`define _INPUT_REPEAT_141 `_INPUT_REPEAT_140 `SET_TEXT_INPUT(140)
`define _INPUT_REPEAT_142 `_INPUT_REPEAT_141 `SET_TEXT_INPUT(141)
`define _INPUT_REPEAT_143 `_INPUT_REPEAT_142 `SET_TEXT_INPUT(142)
`define _INPUT_REPEAT_144 `_INPUT_REPEAT_143 `SET_TEXT_INPUT(143)
`define _INPUT_REPEAT_145 `_INPUT_REPEAT_144 `SET_TEXT_INPUT(144)
`define _INPUT_REPEAT_146 `_INPUT_REPEAT_145 `SET_TEXT_INPUT(145)
`define _INPUT_REPEAT_147 `_INPUT_REPEAT_146 `SET_TEXT_INPUT(146)
`define _INPUT_REPEAT_148 `_INPUT_REPEAT_147 `SET_TEXT_INPUT(147)
`define _INPUT_REPEAT_149 `_INPUT_REPEAT_148 `SET_TEXT_INPUT(148)
`define _INPUT_REPEAT_150 `_INPUT_REPEAT_149 `SET_TEXT_INPUT(149)
`define _INPUT_REPEAT_151 `_INPUT_REPEAT_150 `SET_TEXT_INPUT(150)
`define _INPUT_REPEAT_152 `_INPUT_REPEAT_151 `SET_TEXT_INPUT(151)
`define _INPUT_REPEAT_153 `_INPUT_REPEAT_152 `SET_TEXT_INPUT(152)
`define _INPUT_REPEAT_154 `_INPUT_REPEAT_153 `SET_TEXT_INPUT(153)
`define _INPUT_REPEAT_155 `_INPUT_REPEAT_154 `SET_TEXT_INPUT(154)
`define _INPUT_REPEAT_156 `_INPUT_REPEAT_155 `SET_TEXT_INPUT(155)
`define _INPUT_REPEAT_157 `_INPUT_REPEAT_156 `SET_TEXT_INPUT(156)
`define _INPUT_REPEAT_158 `_INPUT_REPEAT_157 `SET_TEXT_INPUT(157)
`define _INPUT_REPEAT_159 `_INPUT_REPEAT_158 `SET_TEXT_INPUT(158)
`define _INPUT_REPEAT_160 `_INPUT_REPEAT_159 `SET_TEXT_INPUT(159)
`define _INPUT_REPEAT_161 `_INPUT_REPEAT_160 `SET_TEXT_INPUT(160)
`define _INPUT_REPEAT_162 `_INPUT_REPEAT_161 `SET_TEXT_INPUT(161)
`define _INPUT_REPEAT_163 `_INPUT_REPEAT_162 `SET_TEXT_INPUT(162)
`define _INPUT_REPEAT_164 `_INPUT_REPEAT_163 `SET_TEXT_INPUT(163)
`define _INPUT_REPEAT_165 `_INPUT_REPEAT_164 `SET_TEXT_INPUT(164)
`define _INPUT_REPEAT_166 `_INPUT_REPEAT_165 `SET_TEXT_INPUT(165)
`define _INPUT_REPEAT_167 `_INPUT_REPEAT_166 `SET_TEXT_INPUT(166)
`define _INPUT_REPEAT_168 `_INPUT_REPEAT_167 `SET_TEXT_INPUT(167)
`define _INPUT_REPEAT_169 `_INPUT_REPEAT_168 `SET_TEXT_INPUT(168)
`define _INPUT_REPEAT_170 `_INPUT_REPEAT_169 `SET_TEXT_INPUT(169)
`define _INPUT_REPEAT_171 `_INPUT_REPEAT_170 `SET_TEXT_INPUT(170)
`define _INPUT_REPEAT_172 `_INPUT_REPEAT_171 `SET_TEXT_INPUT(171)
`define _INPUT_REPEAT_173 `_INPUT_REPEAT_172 `SET_TEXT_INPUT(172)
`define _INPUT_REPEAT_174 `_INPUT_REPEAT_173 `SET_TEXT_INPUT(173)
`define _INPUT_REPEAT_175 `_INPUT_REPEAT_174 `SET_TEXT_INPUT(174)
`define _INPUT_REPEAT_176 `_INPUT_REPEAT_175 `SET_TEXT_INPUT(175)
`define _INPUT_REPEAT_177 `_INPUT_REPEAT_176 `SET_TEXT_INPUT(176)
`define _INPUT_REPEAT_178 `_INPUT_REPEAT_177 `SET_TEXT_INPUT(177)
`define _INPUT_REPEAT_179 `_INPUT_REPEAT_178 `SET_TEXT_INPUT(178)
`define _INPUT_REPEAT_180 `_INPUT_REPEAT_179 `SET_TEXT_INPUT(179)
`define _INPUT_REPEAT_181 `_INPUT_REPEAT_180 `SET_TEXT_INPUT(180)
`define _INPUT_REPEAT_182 `_INPUT_REPEAT_181 `SET_TEXT_INPUT(181)
`define _INPUT_REPEAT_183 `_INPUT_REPEAT_182 `SET_TEXT_INPUT(182)
`define _INPUT_REPEAT_184 `_INPUT_REPEAT_183 `SET_TEXT_INPUT(183)
`define _INPUT_REPEAT_185 `_INPUT_REPEAT_184 `SET_TEXT_INPUT(184)
`define _INPUT_REPEAT_186 `_INPUT_REPEAT_185 `SET_TEXT_INPUT(185)
`define _INPUT_REPEAT_187 `_INPUT_REPEAT_186 `SET_TEXT_INPUT(186)
`define _INPUT_REPEAT_188 `_INPUT_REPEAT_187 `SET_TEXT_INPUT(187)
`define _INPUT_REPEAT_189 `_INPUT_REPEAT_188 `SET_TEXT_INPUT(188)
`define _INPUT_REPEAT_190 `_INPUT_REPEAT_189 `SET_TEXT_INPUT(189)
`define _INPUT_REPEAT_191 `_INPUT_REPEAT_190 `SET_TEXT_INPUT(190)
`define _INPUT_REPEAT_192 `_INPUT_REPEAT_191 `SET_TEXT_INPUT(191)
`define _INPUT_REPEAT_193 `_INPUT_REPEAT_192 `SET_TEXT_INPUT(192)
`define _INPUT_REPEAT_194 `_INPUT_REPEAT_193 `SET_TEXT_INPUT(193)
`define _INPUT_REPEAT_195 `_INPUT_REPEAT_194 `SET_TEXT_INPUT(194)
`define _INPUT_REPEAT_196 `_INPUT_REPEAT_195 `SET_TEXT_INPUT(195)
`define _INPUT_REPEAT_197 `_INPUT_REPEAT_196 `SET_TEXT_INPUT(196)
`define _INPUT_REPEAT_198 `_INPUT_REPEAT_197 `SET_TEXT_INPUT(197)
`define _INPUT_REPEAT_199 `_INPUT_REPEAT_198 `SET_TEXT_INPUT(198)
`define _INPUT_REPEAT_200 `_INPUT_REPEAT_199 `SET_TEXT_INPUT(199)
`define _INPUT_REPEAT_201 `_INPUT_REPEAT_200 `SET_TEXT_INPUT(200)
`define _INPUT_REPEAT_202 `_INPUT_REPEAT_201 `SET_TEXT_INPUT(201)
`define _INPUT_REPEAT_203 `_INPUT_REPEAT_202 `SET_TEXT_INPUT(202)
`define _INPUT_REPEAT_204 `_INPUT_REPEAT_203 `SET_TEXT_INPUT(203)
`define _INPUT_REPEAT_205 `_INPUT_REPEAT_204 `SET_TEXT_INPUT(204)
`define _INPUT_REPEAT_206 `_INPUT_REPEAT_205 `SET_TEXT_INPUT(205)
`define _INPUT_REPEAT_207 `_INPUT_REPEAT_206 `SET_TEXT_INPUT(206)
`define _INPUT_REPEAT_208 `_INPUT_REPEAT_207 `SET_TEXT_INPUT(207)
`define _INPUT_REPEAT_209 `_INPUT_REPEAT_208 `SET_TEXT_INPUT(208)
`define _INPUT_REPEAT_210 `_INPUT_REPEAT_209 `SET_TEXT_INPUT(209)
`define _INPUT_REPEAT_211 `_INPUT_REPEAT_210 `SET_TEXT_INPUT(210)
`define _INPUT_REPEAT_212 `_INPUT_REPEAT_211 `SET_TEXT_INPUT(211)
`define _INPUT_REPEAT_213 `_INPUT_REPEAT_212 `SET_TEXT_INPUT(212)
`define _INPUT_REPEAT_214 `_INPUT_REPEAT_213 `SET_TEXT_INPUT(213)
`define _INPUT_REPEAT_215 `_INPUT_REPEAT_214 `SET_TEXT_INPUT(214)
`define _INPUT_REPEAT_216 `_INPUT_REPEAT_215 `SET_TEXT_INPUT(215)
`define _INPUT_REPEAT_217 `_INPUT_REPEAT_216 `SET_TEXT_INPUT(216)
`define _INPUT_REPEAT_218 `_INPUT_REPEAT_217 `SET_TEXT_INPUT(217)
`define _INPUT_REPEAT_219 `_INPUT_REPEAT_218 `SET_TEXT_INPUT(218)
`define _INPUT_REPEAT_220 `_INPUT_REPEAT_219 `SET_TEXT_INPUT(219)
`define _INPUT_REPEAT_221 `_INPUT_REPEAT_220 `SET_TEXT_INPUT(220)
`define _INPUT_REPEAT_222 `_INPUT_REPEAT_221 `SET_TEXT_INPUT(221)
`define _INPUT_REPEAT_223 `_INPUT_REPEAT_222 `SET_TEXT_INPUT(222)
`define _INPUT_REPEAT_224 `_INPUT_REPEAT_223 `SET_TEXT_INPUT(223)
`define _INPUT_REPEAT_225 `_INPUT_REPEAT_224 `SET_TEXT_INPUT(224)
`define _INPUT_REPEAT_226 `_INPUT_REPEAT_225 `SET_TEXT_INPUT(225)
`define _INPUT_REPEAT_227 `_INPUT_REPEAT_226 `SET_TEXT_INPUT(226)
`define _INPUT_REPEAT_228 `_INPUT_REPEAT_227 `SET_TEXT_INPUT(227)
`define _INPUT_REPEAT_229 `_INPUT_REPEAT_228 `SET_TEXT_INPUT(228)
`define _INPUT_REPEAT_230 `_INPUT_REPEAT_229 `SET_TEXT_INPUT(229)
`define _INPUT_REPEAT_231 `_INPUT_REPEAT_230 `SET_TEXT_INPUT(230)
`define _INPUT_REPEAT_232 `_INPUT_REPEAT_231 `SET_TEXT_INPUT(231)
`define _INPUT_REPEAT_233 `_INPUT_REPEAT_232 `SET_TEXT_INPUT(232)
`define _INPUT_REPEAT_234 `_INPUT_REPEAT_233 `SET_TEXT_INPUT(233)
`define _INPUT_REPEAT_235 `_INPUT_REPEAT_234 `SET_TEXT_INPUT(234)
`define _INPUT_REPEAT_236 `_INPUT_REPEAT_235 `SET_TEXT_INPUT(235)
`define _INPUT_REPEAT_237 `_INPUT_REPEAT_236 `SET_TEXT_INPUT(236)
`define _INPUT_REPEAT_238 `_INPUT_REPEAT_237 `SET_TEXT_INPUT(237)
`define _INPUT_REPEAT_239 `_INPUT_REPEAT_238 `SET_TEXT_INPUT(238)
`define _INPUT_REPEAT_240 `_INPUT_REPEAT_239 `SET_TEXT_INPUT(239)
`define _INPUT_REPEAT_241 `_INPUT_REPEAT_240 `SET_TEXT_INPUT(240)
`define _INPUT_REPEAT_242 `_INPUT_REPEAT_241 `SET_TEXT_INPUT(241)
`define _INPUT_REPEAT_243 `_INPUT_REPEAT_242 `SET_TEXT_INPUT(242)
`define _INPUT_REPEAT_244 `_INPUT_REPEAT_243 `SET_TEXT_INPUT(243)
`define _INPUT_REPEAT_245 `_INPUT_REPEAT_244 `SET_TEXT_INPUT(244)
`define _INPUT_REPEAT_246 `_INPUT_REPEAT_245 `SET_TEXT_INPUT(245)
`define _INPUT_REPEAT_247 `_INPUT_REPEAT_246 `SET_TEXT_INPUT(246)
`define _INPUT_REPEAT_248 `_INPUT_REPEAT_247 `SET_TEXT_INPUT(247)
`define _INPUT_REPEAT_249 `_INPUT_REPEAT_248 `SET_TEXT_INPUT(248)
`define _INPUT_REPEAT_250 `_INPUT_REPEAT_249 `SET_TEXT_INPUT(249)
`define _INPUT_REPEAT_251 `_INPUT_REPEAT_250 `SET_TEXT_INPUT(250)
`define _INPUT_REPEAT_252 `_INPUT_REPEAT_251 `SET_TEXT_INPUT(251)
`define _INPUT_REPEAT_253 `_INPUT_REPEAT_252 `SET_TEXT_INPUT(252)
`define _INPUT_REPEAT_254 `_INPUT_REPEAT_253 `SET_TEXT_INPUT(253)
`define _INPUT_REPEAT_255 `_INPUT_REPEAT_254 `SET_TEXT_INPUT(254)
`define _INPUT_REPEAT_256 `_INPUT_REPEAT_255 `SET_TEXT_INPUT(255)


`endif